module addr_Writer(
    input wire [9:0] X,
    input wire [9:0] Y,
    input wire [15:0] data,
    input wire [9:0] offset,
    output reg pixelOn
);

    always @(*) begin
              
    end

endmodule
