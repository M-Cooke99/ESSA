module Test()

end module